module BloodyRoot ();

	DataPath dp (.(*));
	ControlPath cp (.(*));

endmodule : BloodyRoot