module system_tb();


endmodule : system_tb