module ControlPath();

endmodule : ControlPath