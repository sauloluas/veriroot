module Top ();

	BloodyRoot br (.(*));
	Ram dmem (.(*));
	Rom imem (.(*));


endmodule : Top